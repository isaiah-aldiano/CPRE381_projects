-------------------------------------------------------------------------
-- Sam Burns 
-- Department of Electrical and Computer Engineering
-- Iowa State University
-------------------------------------------------------------------------


-- Decoder5to32.vhd
-------------------------------------------------------------------------
-- DESCRIPTION: This file contains an implementation of a 5 to 32 decoder 
-- using "with-select" statements
--
--
-- NOTES:
-- created 17:15 2/6/2025
-------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity Decoder5to32 is 
   port(sel : in std_logic_vector(4 downto 0);
      write_en : in std_logic;
   	out_sel : out std_logic_vector(31 downto 0));
end Decoder5to32;

architecture behavioral of Decoder5to32 is 

   signal p1_out : std_logic_vector(31 downto 0);
   begin 
--Use with select statements for 5 bit input to 32 bit output assignment
   with sel select
      p1_out <=   "00000000000000000000000000000001" when "00000",
                   "00000000000000000000000000000010" when "00001",
                   "00000000000000000000000000000100" when "00010",
                   "00000000000000000000000000001000" when "00011",
                   "00000000000000000000000000010000" when "00100",
                   "00000000000000000000000000100000" when "00101",
                   "00000000000000000000000001000000" when "00110",
                   "00000000000000000000000010000000" when "00111",
                   "00000000000000000000000100000000" when "01000",
                   "00000000000000000000001000000000" when "01001",
                   "00000000000000000000010000000000" when "01010",
                   "00000000000000000000100000000000" when "01011",
                   "00000000000000000001000000000000" when "01100",
                   "00000000000000000010000000000000" when "01101",
                   "00000000000000000100000000000000" when "01110",
                   "00000000000000001000000000000000" when "01111",
                   "00000000000000010000000000000000" when "10000",
                   "00000000000000100000000000000000" when "10001",
                   "00000000000001000000000000000000" when "10010",
                   "00000000000010000000000000000000" when "10011",
                   "00000000000100000000000000000000" when "10100",
                   "00000000001000000000000000000000" when "10101",
                   "00000000010000000000000000000000" when "10110",
                   "00000000100000000000000000000000" when "10111",
                   "00000001000000000000000000000000" when "11000",
                   "00000010000000000000000000000000" when "11001",
                   "00000100000000000000000000000000" when "11010",
                   "00001000000000000000000000000000" when "11011",
                   "00010000000000000000000000000000" when "11100",
                   "00100000000000000000000000000000" when "11101",
                   "01000000000000000000000000000000" when "11110",
                   "10000000000000000000000000000000" when "11111",
                   (others => '0') when others; -- Default case

   with write_en select
      out_sel <= "00000000000000000000000000000000" when '0',
                 p1_out when '1',
                 (others => '0') when others;

   
end behavioral;
